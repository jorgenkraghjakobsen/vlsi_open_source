module top(input [2:0] op0, input [2:0] op1, output [5:0] result);
    assign result = op0 * op1;
endmodule
